module dm 
(
  // Declarar os pinos de IO
);

endmodule