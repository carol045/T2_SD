module top 
(
  // Declarar os pinos de IO
);

endmodule