module wrapper 
(
  // Declarar os pinos de IO
);

endmodule