module fibonacci 
(
  // Declarar os pinos de IO
);

endmodule